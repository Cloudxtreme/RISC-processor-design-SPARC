/**************************************
* Module: RegisterWindow
* Date:2014-09-27  
* Author: josediaz     
*
* Description: Register window module
***************************************/
module  RegisterWindow();


endmodule

